`timescale 1ns / 1ps

module instr_decoder( 
    input [31:0] inst,
    output reg [31:0] choose
    );
    always @(*) 
    begin
    if(inst[31:26] == 6'b0)begin
        if(inst[5:0] == 6'b100000)     choose = 32'b0000_0000_0000_0000_0000_0000_0000_0001;//add
        else if(inst[5:0] == 6'b100001)choose = 32'b0000_0000_0000_0000_0000_0000_0000_0010;//addu
        else if(inst[5:0] == 6'b100010)choose = 32'b0000_0000_0000_0000_0000_0000_0000_0100;//sub
        else if(inst[5:0] == 6'b100011)choose = 32'b0000_0000_0000_0000_0000_0000_0000_1000;//subu
        else if(inst[5:0] == 6'b100100)choose = 32'b0000_0000_0000_0000_0000_0000_0001_0000;//and
        else if(inst[5:0] == 6'b100101)choose = 32'b0000_0000_0000_0000_0000_0000_0010_0000;//or
        else if(inst[5:0] == 6'b100110)choose = 32'b0000_0000_0000_0000_0000_0000_0100_0000;//xor
        else if(inst[5:0] == 6'b100111)choose = 32'b0000_0000_0000_0000_0000_0000_1000_0000;//nor
        else if(inst[5:0] == 6'b101010)choose = 32'b0000_0000_0000_0000_0000_0001_0000_0000;//slt
        else if(inst[5:0] == 6'b101011)choose = 32'b0000_0000_0000_0000_0000_0010_0000_0000;//sltu
        else if(inst[5:0] == 6'b000000)choose = 32'b0000_0000_0000_0000_0000_0100_0000_0000;//sll
        else if(inst[5:0] == 6'b000010)choose = 32'b0000_0000_0000_0000_0000_1000_0000_0000;//srl
        else if(inst[5:0] == 6'b000011)choose = 32'b0000_0000_0000_0000_0001_0000_0000_0000;//sra
        else if(inst[5:0] == 6'b000100)choose = 32'b0000_0000_0000_0000_0010_0000_0000_0000;//sllv
        else if(inst[5:0] == 6'b000110)choose = 32'b0000_0000_0000_0000_0100_0000_0000_0000;//srlv
        else if(inst[5:0] == 6'b000111)choose = 32'b0000_0000_0000_0000_1000_0000_0000_0000;//srav
        else if(inst[5:0] == 6'b001000)choose = 32'b0000_0000_0000_0001_0000_0000_0000_0000;//jr
    end
    else if(inst[31:26] == 6'b001000)choose = 32'b0000_0000_0000_0010_0000_0000_0000_0000;//addi
    else if(inst[31:26] == 6'b001001)choose = 32'b0000_0000_0000_0100_0000_0000_0000_0000;//addiu
    else if(inst[31:26] == 6'b001100)choose = 32'b0000_0000_0000_1000_0000_0000_0000_0000;//andi
    else if(inst[31:26] == 6'b001101)choose = 32'b0000_0000_0001_0000_0000_0000_0000_0000;//ori
    else if(inst[31:26] == 6'b001110)choose = 32'b0000_0000_0010_0000_0000_0000_0000_0000;//xori
    else if(inst[31:26] == 6'b100011)choose = 32'b0000_0000_0100_0000_0000_0000_0000_0000;//lw
    else if(inst[31:26] == 6'b101011)choose = 32'b0000_0000_1000_0000_0000_0000_0000_0000;//sw
    else if(inst[31:26] == 6'b000100)choose = 32'b0000_0001_0000_0000_0000_0000_0000_0000;//beq
    else if(inst[31:26] == 6'b000101)choose = 32'b0000_0010_0000_0000_0000_0000_0000_0000;//bne
    else if(inst[31:26] == 6'b001010)choose = 32'b0000_0100_0000_0000_0000_0000_0000_0000;//slti
    else if(inst[31:26] == 6'b001011)choose = 32'b0000_1000_0000_0000_0000_0000_0000_0000;//sltiu
    else if(inst[31:26] == 6'b001111)choose = 32'b0001_0000_0000_0000_0000_0000_0000_0000;//lui
    else if(inst[31:26] == 6'b000010)choose = 32'b0010_0000_0000_0000_0000_0000_0000_0000;//j
    else if(inst[31:26] == 6'b000011)choose = 32'b0100_0000_0000_0000_0000_0000_0000_0000;//jal
    else choose = 32'bz;
    end

endmodule
